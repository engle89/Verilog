`timescale 1ns / 1ps

module ALU2_tb();

	reg [15:0] A, B;
	reg [3:0] ALU_Control;
	
	wire Overflow, Zero;
	wire [15:0] S;
	
	ALU2 uut(A, B, ALU_Control, Overflow, Zero, S);
	
	initial begin
		A = 0;
		B = 0;
		ALU_Control = 0;
		
		// Subtraction
		#10 ALU_Control = 4'b0000;
		A = 	  16'b0000000000000001; B=16'b0000000000000001;	// 0
		#10 A = 16'b0000000000000010; B=16'b0000000000000001;	// 1
		#10 A = 16'b0000000000000000; B=16'b0000000000000001;	// all 1s
		#10 A = 16'b1000000000000000; B=16'b0111111111111111;
		
		// Addition
		#10 ALU_Control = 4'b0001;
		A =     16'b0000000000000001; B=16'b0000000000000001;		// 10
		#10 A = 16'b0000000000000001; B=16'b0000000000000010;	// 11
		#10 A = 16'b1111111111111111; B=16'b0000000000000001;	// all 0s, overflow 1
		#10 A = 16'b0111111111111111; B=16'b0000000000000001;
		
		// Bitwise Or
		#10 ALU_Control = 4'b0010;
		A =     16'b0000000000000001; B=16'b0000000000000001;		// 1
		#10 A = 16'b0000000000000001; B=16'b0000000000000010;	// 11
		#10 A = 16'b1111111111111111; B=16'b0000000000000001; // all 1s
		
		// Bitwise And
		#10 ALU_Control = 4'b0011;
		A =     16'b0000000000000001; B=16'b0000000000000001;		// 1
		#10 A = 16'b0000000000000001; B=16'b0000000000000100;	// all 0s
		#10 A = 16'b1111111111111111; B=16'b0000000000000001; // 1
		
		// Decrement
		#10 ALU_Control = 4'b0100;
		A =     16'b0000000000000001; B=16'b0000000000000001;		// 0
		#10 A = 16'b0000000000000000; B=16'b0000000000000001;	// all 1s
		#10 A=  16'b1000000000000000;
		
		// Increment
		#10 ALU_Control = 4'b0101;
		A =     16'b0000000000000001; B=16'b0000000000000010;	// 10
		#10 A = 16'b0111111111111111; B=16'b0000000000000001;	// 1 with 15 0s
		#10 A = 16'b1111111111111111; B=16'b0000000000000001;	// all 0s, overflow 1
		
		// Invert
		#10 ALU_Control = 4'b0110;
		A =     16'b0000000000000001; B=16'b000000000000010;
		#10 A = 16'b0111111111111111; B=16'b0000000000000001;
		
		// Arithmetic Left Shift
		#10 ALU_Control = 4'b1100;
		A =     16'b0000000000000001; B=16'b0000000000000010;	// 100
		#10 A = 16'b0111111111111111; B=16'b0000000000000001;
		#10 A = 16'b1111111111111111; B=16'b0000000000000001;
		
		// Arithmetic Right Shift
		#10 ALU_Control = 4'b1110;
		A =     16'b0000000000000010; B=16'b0000000000000001;	// 1
		#10 A = 16'b0111111111111111; B=16'b0000000000000001;
		#10 A = 16'b1111111111111111; B=16'b0000000000000001;
		
		// Logical Left Shift
		#10 ALU_Control = 4'b1000;
		A =     16'b0000000000000001; B=16'b0000000000000010;	// 100
		#10 A = 16'b0111111111111111; B=16'b0000000000000001;
		#10 A = 16'b1111111111111111; B=16'b0000000000000001;
		
		// Logical Right Shift
		#10 ALU_Control = 4'b1010;
		A =     16'b0000000000000010; B=16'b0000000000000001;
		#10 A = 16'b0111111111111111; B=16'b0000000000000001;
		#10 A = 16'b1111111111111111; B=16'b0000000000000001;
		
		// Set On Less Than or Equal
		#10 ALU_Control = 4'b1001;
		A =     16'b0000000000000010; B=16'b0000000000000001; // 0
		#10 A = 16'b0000000000000010; B=16'b0000000000000100;	// 1
		#10 A = 16'b1111111111111111; B=16'b1111111111111111; // 1
		#10 A = 16'b0111111111111111; B=16'b1111111111111111;
		
	end

endmodule
